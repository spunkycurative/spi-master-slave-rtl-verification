class driver;
  
  // Virtual interface handle to connect to the DUT's pins
  virtual spi_if vif;
  
  // Local transaction object (will hold the transaction fetched from the generator)
  transaction tr;
  
  // Mailbox to get the transaction objects from the generator
  mailbox #(transaction) mbx;
  
  // Mailbox to send the expected DIN (Data In) to the scoreboard/checker
  // The Data Structure (DS) is a simple 12-bit value in this case.
  mailbox #(bit [11:0]) mbxds;
  
  // Event: Signal for flow control (currently unused, but good for complex control)
  event drvnext;
  
  // A local variable to hold data if needed (currently unused, but kept for clarity)
  bit [11:0] din;
  
  // Constructor: Initializes the mailboxes
  function new (mailbox #(bit [11:0]) mbxds, mailbox #(transaction) mbx);
    this.mbx = mbx;
    this.mbxds = mbxds;
  endfunction
  
  // Task to handle the active-low reset sequence
  task reset();
    // 1. Assert reset and initialize interface signals to a known state
    vif.rst <= 1'b1;
    vif.newd <= 1'b0;
    vif.din <= 1'b0;
    
    // 2. Hold reset for 10 clock cycles
    repeat(10) @(posedge vif.clk);
    
    // 3. De-assert reset
    vif.rst <= 1'b0;
    
    // 4. Wait for 5 more clock cycles for system stabilization
    repeat(5) @(posedge vif.clk);
    
  endtask
  
  // Main task to drive transactions
  task run();
    
    forever begin
      // 1. Get a new randomized transaction from the generator's mailbox
      mbx.get(tr);
      
      // 2. Wait for the SPI clock edge (assuming SCLK is generated by the master)
      @(posedge vif.sclk);
      
      // 3. Drive the stimulus: Assert newd and put the data onto the din bus
      vif.newd <= 1'b1;
      vif.din <= tr.din;
      
      // 4. Send the expected input data to the scoreboard
      // This is crucial: the scoreboard needs the *input* to predict the *output*.
      mbxds.put(tr.din);
      
      // 5. Wait for the next SCLK edge to de-assert newd
      @(posedge vif.sclk);
      vif.newd <= 1'b0;
      
      // 6. Wait for the DUT's done signal to confirm the transfer is complete
      @(posedge vif.done);
      
      $display("[DRV]: data sent to DUT = %0d", tr.din);
      
      // 7. Wait one more SCLK cycle before looking for the next transaction
      @(posedge vif.sclk);
      
    end
  endtask
  
endclass
